module imem #(parameter N = 32)(
    input logic[7:0] addr0, addr1,
    output logic[N-1:0] q0, q1
);
    logic [N - 1:0] rom [0 : 255];
    assign rom[0:145] = '{
        32'h00003197, //   0: auipc gp,0x3
        32'h00018193, //   4: mv gp,gp
        32'h00003023, //   8: sd zero,0(zero) # 0 <start>
        32'h00002117, //   c: auipc sp,0x2
        32'hff410113, //  10: addi sp,sp,-12 # 2000 <stack_top>
        32'h00010413, //  14: mv s0,sp
        32'h00010fb7, //  18: lui t6,0x10
        32'hff8f8f9b, //  1c: addiw t6,t6,-8 # fff8 <global_pointer+0xcff8>
        32'h000fbf03, //  20: ld t5,0(t6)
        32'h00018493, //  24: mv s1,gp
        32'hff0f8f93, //  28: addi t6,t6,-16
        32'h00848493, //  2c: addi s1,s1,8
        32'h000fbe83, //  30: ld t4,0(t6)
        32'h008fbe03, //  34: ld t3,8(t6)
        32'h020e9e93, //  38: slli t4,t4,0x20
        32'h01de0e33, //  3c: add t3,t3,t4
        32'h01c4b023, //  40: sd t3,0(s1)
        32'hffff0f13, //  44: addi t5,t5,-1
        32'hfe0f10e3, //  48: bnez t5,28 <rom_read>
        32'h30046073, //  4c: csrsi mstatus,8
        32'h00000f17, //  50: auipc t5,0x0
        32'h01cf0f13, //  54: addi t5,t5,28 # 6c <never_ret>
        32'h305f1073, //  58: csrw mtvec,t5
        32'h154000ef, //  5c: jal ra,1b0 <main>
        32'h00100f93, //  60: li t6,1
        32'h01f03023, //  64: sd t6,0(zero) # 0 <start>
        32'h00100073, //  68: ebreak
        32'h0000006f, //  6c: j 6c <never_ret>
        32'hfc010113, //  70: addi sp,sp,-64
        32'h02813c23, //  74: sd s0,56(sp)
        32'h00000013, //  78: nop
        32'h04010413, //  7c: addi s0,sp,64
        32'hfca43c23, //  80: sd a0,-40(s0)
        32'h00000013, //  84: nop
        32'hfcb43823, //  88: sd a1,-48(s0)
        32'h00000013, //  8c: nop
        32'h00060793, //  90: mv a5,a2
        32'hfcf42623, //  94: sw a5,-52(s0)
        32'hfd843783, //  98: ld a5,-40(s0)
        32'hfd843783, //  9c: ld a5,-40(s0)
        32'hfef43423, //  a0: sd a5,-24(s0)
        32'h00000013, //  a4: nop
        32'hfd043783, //  a8: ld a5,-48(s0)
        32'hfd043783, //  ac: ld a5,-48(s0)
        32'hfef43023, //  b0: sd a5,-32(s0)
        32'h00000013, //  b4: nop
        32'h0400006f, //  b8: j f8 <memcpy+0x88>
        32'hfe043703, //  bc: ld a4,-32(s0)
        32'hfe043703, //  c0: ld a4,-32(s0)
        32'h00170793, //  c4: addi a5,a4,1
        32'hfef43023, //  c8: sd a5,-32(s0)
        32'h00000013, //  cc: nop
        32'hfe843783, //  d0: ld a5,-24(s0)
        32'hfe843783, //  d4: ld a5,-24(s0)
        32'h00178693, //  d8: addi a3,a5,1
        32'hfed43423, //  dc: sd a3,-24(s0)
        32'h00000013, //  e0: nop
        32'h00074703, //  e4: lbu a4,0(a4)
        32'h00e78023, //  e8: sb a4,0(a5)
        32'hfcc42783, //  ec: lw a5,-52(s0)
        32'hfff7879b, //  f0: addiw a5,a5,-1
        32'hfcf42623, //  f4: sw a5,-52(s0)
        32'hfcc42783, //  f8: lw a5,-52(s0)
        32'h0007879b, //  fc: sext.w a5,a5
        32'hfa079ee3, // 100: bnez a5,bc <memcpy+0x4c>
        32'hfd843783, // 104: ld a5,-40(s0)
        32'hfd843783, // 108: ld a5,-40(s0)
        32'h00078513, // 10c: mv a0,a5
        32'h03813403, // 110: ld s0,56(sp)
        32'h03813403, // 114: ld s0,56(sp)
        32'h04010113, // 118: addi sp,sp,64
        32'h00008067, // 11c: ret
        32'hfd010113, // 120: addi sp,sp,-48
        32'h02813423, // 124: sd s0,40(sp)
        32'h00000013, // 128: nop
        32'h03010413, // 12c: addi s0,sp,48
        32'hfca43c23, // 130: sd a0,-40(s0)
        32'h00000013, // 134: nop
        32'hfe043423, // 138: sd zero,-24(s0)
        32'h00000013, // 13c: nop
        32'h00100793, // 140: li a5,1
        32'hfef43023, // 144: sd a5,-32(s0)
        32'h00000013, // 148: nop
        32'h0340006f, // 14c: j 180 <sum+0x60>
        32'hfe843703, // 150: ld a4,-24(s0)
        32'hfe843703, // 154: ld a4,-24(s0)
        32'hfe043783, // 158: ld a5,-32(s0)
        32'hfe043783, // 15c: ld a5,-32(s0)
        32'h00f707b3, // 160: add a5,a4,a5
        32'hfef43423, // 164: sd a5,-24(s0)
        32'h00000013, // 168: nop
        32'hfe043783, // 16c: ld a5,-32(s0)
        32'hfe043783, // 170: ld a5,-32(s0)
        32'h00178793, // 174: addi a5,a5,1
        32'hfef43023, // 178: sd a5,-32(s0)
        32'h00000013, // 17c: nop
        32'hfe043703, // 180: ld a4,-32(s0)
        32'hfe043703, // 184: ld a4,-32(s0)
        32'hfd843783, // 188: ld a5,-40(s0)
        32'hfd843783, // 18c: ld a5,-40(s0)
        32'hfce7f0e3, // 190: bgeu a5,a4,150 <sum+0x30>
        32'hfe843783, // 194: ld a5,-24(s0)
        32'hfe843783, // 198: ld a5,-24(s0)
        32'h00078513, // 19c: mv a0,a5
        32'h02813403, // 1a0: ld s0,40(sp)
        32'h02813403, // 1a4: ld s0,40(sp)
        32'h03010113, // 1a8: addi sp,sp,48
        32'h00008067, // 1ac: ret
        32'hf4010113, // 1b0: addi sp,sp,-192
        32'h0a113c23, // 1b4: sd ra,184(sp)
        32'h00000013, // 1b8: nop
        32'h0a813823, // 1bc: sd s0,176(sp)
        32'h00000013, // 1c0: nop
        32'h0c010413, // 1c4: addi s0,sp,192
        32'h000037b7, // 1c8: lui a5,0x3
        32'h00078713, // 1cc: mv a4,a5
        32'hf4840793, // 1d0: addi a5,s0,-184
        32'h00070693, // 1d4: mv a3,a4
        32'h09800713, // 1d8: li a4,152
        32'h00070613, // 1dc: mv a2,a4
        32'h00068593, // 1e0: mv a1,a3
        32'h00078513, // 1e4: mv a0,a5
        32'he89ff0ef, // 1e8: jal ra,70 <memcpy>
        32'h00000013, // 1ec: nop
        32'h00000013, // 1f0: nop
        32'h00000013, // 1f4: nop
        32'hf4843783, // 1f8: ld a5,-184(s0)
        32'hf4843783, // 1fc: ld a5,-184(s0)
        32'hfef43423, // 200: sd a5,-24(s0)
        32'h00000013, // 204: nop
        32'h00000013, // 208: nop
        32'h00000013, // 20c: nop
        32'h00000013, // 210: nop
        32'h00a00513, // 214: li a0,10
        32'hf09ff0ef, // 218: jal ra,120 <sum>
        32'hfea43023, // 21c: sd a0,-32(s0)
        32'h00000013, // 220: nop
        32'hfe043783, // 224: ld a5,-32(s0)
        32'hfe043783, // 228: ld a5,-32(s0)
        32'h00078513, // 22c: mv a0,a5
        32'h0b813083, // 230: ld ra,184(sp)
        32'h0b813083, // 234: ld ra,184(sp)
        32'h0b013403, // 238: ld s0,176(sp)
        32'h0b013403, // 23c: ld s0,176(sp)
        32'h0c010113, // 240: addi sp,sp,192
        32'h00008067 // 244: ret
    };
    assign rom[217:255] = '{
        32'h00000000,
        32'h00000006,
        32'h00000000,
        32'h00000005,
        32'h00000000,
        32'h00000002,
        32'h00000000,
        32'h00000001,
        32'h00000000,
        32'h00000005,
        32'h00000000,
        32'h0000007b,
        32'h00000000,
        32'h000001b0,
        32'h00000000,
        32'h00000002,
        32'h00000000,
        32'h00000001,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000009,
        32'h00000000,
        32'h00000008,
        32'h00000000,
        32'h00000007,
        32'h00000000,
        32'h00000006,
        32'h00000000,
        32'h00000005,
        32'h00000000,
        32'h00000004,
        32'h00000000,
        32'h00000003,
        32'h00000000,
        32'h00000002,
        32'h00000001,
        32'h00000007,
        32'h13
    };
    assign rom [146:216] = '{(71){'0}};
    assign q0 = rom[addr0];
    assign q1 = rom[addr1];
endmodule