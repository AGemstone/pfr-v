// coprocessor.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module coprocessor (
		input  wire        clk_clk,                //             clk.clk
		output wire [14:0] pio_addr_export,        //        pio_addr.export
		output wire [5:0]  pio_control_export,     //     pio_control.export
		input  wire [31:0] pio_data_high_in_port,  //   pio_data_high.in_port
		output wire [31:0] pio_data_high_out_port, //                .out_port
		input  wire [31:0] pio_data_low_in_port,   //    pio_data_low.in_port
		output wire [31:0] pio_data_low_out_port,  //                .out_port
		input  wire [1:0]  pio_riscv_flags_export, // pio_riscv_flags.export
		input  wire        reset_reset_n           //           reset.reset_n
	);

	wire  [31:0] niosii_data_master_readdata;                               // mm_interconnect_0:NiosII_data_master_readdata -> NiosII:d_readdata
	wire         niosii_data_master_waitrequest;                            // mm_interconnect_0:NiosII_data_master_waitrequest -> NiosII:d_waitrequest
	wire         niosii_data_master_debugaccess;                            // NiosII:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NiosII_data_master_debugaccess
	wire  [14:0] niosii_data_master_address;                                // NiosII:d_address -> mm_interconnect_0:NiosII_data_master_address
	wire   [3:0] niosii_data_master_byteenable;                             // NiosII:d_byteenable -> mm_interconnect_0:NiosII_data_master_byteenable
	wire         niosii_data_master_read;                                   // NiosII:d_read -> mm_interconnect_0:NiosII_data_master_read
	wire         niosii_data_master_write;                                  // NiosII:d_write -> mm_interconnect_0:NiosII_data_master_write
	wire  [31:0] niosii_data_master_writedata;                              // NiosII:d_writedata -> mm_interconnect_0:NiosII_data_master_writedata
	wire  [31:0] niosii_instruction_master_readdata;                        // mm_interconnect_0:NiosII_instruction_master_readdata -> NiosII:i_readdata
	wire         niosii_instruction_master_waitrequest;                     // mm_interconnect_0:NiosII_instruction_master_waitrequest -> NiosII:i_waitrequest
	wire  [14:0] niosii_instruction_master_address;                         // NiosII:i_address -> mm_interconnect_0:NiosII_instruction_master_address
	wire         niosii_instruction_master_read;                            // NiosII:i_read -> mm_interconnect_0:NiosII_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_readdata;         // NiosII:debug_mem_slave_readdata -> mm_interconnect_0:NiosII_debug_mem_slave_readdata
	wire         mm_interconnect_0_niosii_debug_mem_slave_waitrequest;      // NiosII:debug_mem_slave_waitrequest -> mm_interconnect_0:NiosII_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_niosii_debug_mem_slave_debugaccess;      // mm_interconnect_0:NiosII_debug_mem_slave_debugaccess -> NiosII:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_niosii_debug_mem_slave_address;          // mm_interconnect_0:NiosII_debug_mem_slave_address -> NiosII:debug_mem_slave_address
	wire         mm_interconnect_0_niosii_debug_mem_slave_read;             // mm_interconnect_0:NiosII_debug_mem_slave_read -> NiosII:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_niosii_debug_mem_slave_byteenable;       // mm_interconnect_0:NiosII_debug_mem_slave_byteenable -> NiosII:debug_mem_slave_byteenable
	wire         mm_interconnect_0_niosii_debug_mem_slave_write;            // mm_interconnect_0:NiosII_debug_mem_slave_write -> NiosII:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_writedata;        // mm_interconnect_0:NiosII_debug_mem_slave_writedata -> NiosII:debug_mem_slave_writedata
	wire         mm_interconnect_0_memory_s1_chipselect;                    // mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                      // memory:readdata -> mm_interconnect_0:memory_s1_readdata
	wire  [10:0] mm_interconnect_0_memory_s1_address;                       // mm_interconnect_0:memory_s1_address -> memory:address
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;                    // mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	wire         mm_interconnect_0_memory_s1_write;                         // mm_interconnect_0:memory_s1_write -> memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                     // mm_interconnect_0:memory_s1_writedata -> memory:writedata
	wire         mm_interconnect_0_memory_s1_clken;                         // mm_interconnect_0:memory_s1_clken -> memory:clken
	wire         mm_interconnect_0_io_data_low_s1_chipselect;               // mm_interconnect_0:io_data_low_s1_chipselect -> io_data_low:chipselect
	wire  [31:0] mm_interconnect_0_io_data_low_s1_readdata;                 // io_data_low:readdata -> mm_interconnect_0:io_data_low_s1_readdata
	wire   [1:0] mm_interconnect_0_io_data_low_s1_address;                  // mm_interconnect_0:io_data_low_s1_address -> io_data_low:address
	wire         mm_interconnect_0_io_data_low_s1_write;                    // mm_interconnect_0:io_data_low_s1_write -> io_data_low:write_n
	wire  [31:0] mm_interconnect_0_io_data_low_s1_writedata;                // mm_interconnect_0:io_data_low_s1_writedata -> io_data_low:writedata
	wire         mm_interconnect_0_io_data_high_s1_chipselect;              // mm_interconnect_0:io_data_high_s1_chipselect -> io_data_high:chipselect
	wire  [31:0] mm_interconnect_0_io_data_high_s1_readdata;                // io_data_high:readdata -> mm_interconnect_0:io_data_high_s1_readdata
	wire   [1:0] mm_interconnect_0_io_data_high_s1_address;                 // mm_interconnect_0:io_data_high_s1_address -> io_data_high:address
	wire         mm_interconnect_0_io_data_high_s1_write;                   // mm_interconnect_0:io_data_high_s1_write -> io_data_high:write_n
	wire  [31:0] mm_interconnect_0_io_data_high_s1_writedata;               // mm_interconnect_0:io_data_high_s1_writedata -> io_data_high:writedata
	wire         mm_interconnect_0_io_addr_s1_chipselect;                   // mm_interconnect_0:io_addr_s1_chipselect -> io_addr:chipselect
	wire  [31:0] mm_interconnect_0_io_addr_s1_readdata;                     // io_addr:readdata -> mm_interconnect_0:io_addr_s1_readdata
	wire   [1:0] mm_interconnect_0_io_addr_s1_address;                      // mm_interconnect_0:io_addr_s1_address -> io_addr:address
	wire         mm_interconnect_0_io_addr_s1_write;                        // mm_interconnect_0:io_addr_s1_write -> io_addr:write_n
	wire  [31:0] mm_interconnect_0_io_addr_s1_writedata;                    // mm_interconnect_0:io_addr_s1_writedata -> io_addr:writedata
	wire         mm_interconnect_0_io_control_s1_chipselect;                // mm_interconnect_0:io_control_s1_chipselect -> io_control:chipselect
	wire  [31:0] mm_interconnect_0_io_control_s1_readdata;                  // io_control:readdata -> mm_interconnect_0:io_control_s1_readdata
	wire   [1:0] mm_interconnect_0_io_control_s1_address;                   // mm_interconnect_0:io_control_s1_address -> io_control:address
	wire         mm_interconnect_0_io_control_s1_write;                     // mm_interconnect_0:io_control_s1_write -> io_control:write_n
	wire  [31:0] mm_interconnect_0_io_control_s1_writedata;                 // mm_interconnect_0:io_control_s1_writedata -> io_control:writedata
	wire  [31:0] mm_interconnect_0_io_riscv_flags_s1_readdata;              // io_riscv_flags:readdata -> mm_interconnect_0:io_riscv_flags_s1_readdata
	wire   [1:0] mm_interconnect_0_io_riscv_flags_s1_address;               // mm_interconnect_0:io_riscv_flags_s1_address -> io_riscv_flags:address
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] niosii_irq_irq;                                            // irq_mapper:sender_irq -> NiosII:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [NiosII:reset_n, io_addr:reset_n, io_control:reset_n, io_data_high:reset_n, io_data_low:reset_n, io_riscv_flags:reset_n, irq_mapper:reset, jtag_uart:rst_n, memory:reset, mm_interconnect_0:NiosII_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [NiosII:reset_req, memory:reset_req, rst_translator:reset_req_in]
	wire         niosii_debug_reset_request_reset;                          // NiosII:debug_reset_request -> rst_controller:reset_in1

	coprocessor_NiosII niosii (
		.clk                                 (clk_clk),                                              //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (niosii_data_master_address),                           //               data_master.address
		.d_byteenable                        (niosii_data_master_byteenable),                        //                          .byteenable
		.d_read                              (niosii_data_master_read),                              //                          .read
		.d_readdata                          (niosii_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (niosii_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (niosii_data_master_write),                             //                          .write
		.d_writedata                         (niosii_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (niosii_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (niosii_instruction_master_address),                    //        instruction_master.address
		.i_read                              (niosii_instruction_master_read),                       //                          .read
		.i_readdata                          (niosii_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (niosii_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (niosii_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (niosii_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_niosii_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_niosii_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_niosii_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_niosii_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_niosii_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_niosii_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_niosii_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_niosii_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	coprocessor_io_addr io_addr (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_io_addr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_io_addr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_io_addr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_io_addr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_io_addr_s1_readdata),   //                    .readdata
		.out_port   (pio_addr_export)                          // external_connection.export
	);

	coprocessor_io_control io_control (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_io_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_io_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_io_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_io_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_io_control_s1_readdata),   //                    .readdata
		.out_port   (pio_control_export)                          // external_connection.export
	);

	coprocessor_io_data_high io_data_high (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_io_data_high_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_io_data_high_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_io_data_high_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_io_data_high_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_io_data_high_s1_readdata),   //                    .readdata
		.in_port    (pio_data_high_in_port),                        // external_connection.export
		.out_port   (pio_data_high_out_port)                        //                    .export
	);

	coprocessor_io_data_high io_data_low (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_io_data_low_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_io_data_low_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_io_data_low_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_io_data_low_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_io_data_low_s1_readdata),   //                    .readdata
		.in_port    (pio_data_low_in_port),                        // external_connection.export
		.out_port   (pio_data_low_out_port)                        //                    .export
	);

	coprocessor_io_riscv_flags io_riscv_flags (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_io_riscv_flags_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_io_riscv_flags_s1_readdata), //                    .readdata
		.in_port  (pio_riscv_flags_export)                        // external_connection.export
	);

	coprocessor_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	coprocessor_memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	coprocessor_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                            (clk_clk),                                                   //                          clk_0_clk.clk
		.NiosII_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // NiosII_reset_reset_bridge_in_reset.reset
		.NiosII_data_master_address               (niosii_data_master_address),                                //                 NiosII_data_master.address
		.NiosII_data_master_waitrequest           (niosii_data_master_waitrequest),                            //                                   .waitrequest
		.NiosII_data_master_byteenable            (niosii_data_master_byteenable),                             //                                   .byteenable
		.NiosII_data_master_read                  (niosii_data_master_read),                                   //                                   .read
		.NiosII_data_master_readdata              (niosii_data_master_readdata),                               //                                   .readdata
		.NiosII_data_master_write                 (niosii_data_master_write),                                  //                                   .write
		.NiosII_data_master_writedata             (niosii_data_master_writedata),                              //                                   .writedata
		.NiosII_data_master_debugaccess           (niosii_data_master_debugaccess),                            //                                   .debugaccess
		.NiosII_instruction_master_address        (niosii_instruction_master_address),                         //          NiosII_instruction_master.address
		.NiosII_instruction_master_waitrequest    (niosii_instruction_master_waitrequest),                     //                                   .waitrequest
		.NiosII_instruction_master_read           (niosii_instruction_master_read),                            //                                   .read
		.NiosII_instruction_master_readdata       (niosii_instruction_master_readdata),                        //                                   .readdata
		.io_addr_s1_address                       (mm_interconnect_0_io_addr_s1_address),                      //                         io_addr_s1.address
		.io_addr_s1_write                         (mm_interconnect_0_io_addr_s1_write),                        //                                   .write
		.io_addr_s1_readdata                      (mm_interconnect_0_io_addr_s1_readdata),                     //                                   .readdata
		.io_addr_s1_writedata                     (mm_interconnect_0_io_addr_s1_writedata),                    //                                   .writedata
		.io_addr_s1_chipselect                    (mm_interconnect_0_io_addr_s1_chipselect),                   //                                   .chipselect
		.io_control_s1_address                    (mm_interconnect_0_io_control_s1_address),                   //                      io_control_s1.address
		.io_control_s1_write                      (mm_interconnect_0_io_control_s1_write),                     //                                   .write
		.io_control_s1_readdata                   (mm_interconnect_0_io_control_s1_readdata),                  //                                   .readdata
		.io_control_s1_writedata                  (mm_interconnect_0_io_control_s1_writedata),                 //                                   .writedata
		.io_control_s1_chipselect                 (mm_interconnect_0_io_control_s1_chipselect),                //                                   .chipselect
		.io_data_high_s1_address                  (mm_interconnect_0_io_data_high_s1_address),                 //                    io_data_high_s1.address
		.io_data_high_s1_write                    (mm_interconnect_0_io_data_high_s1_write),                   //                                   .write
		.io_data_high_s1_readdata                 (mm_interconnect_0_io_data_high_s1_readdata),                //                                   .readdata
		.io_data_high_s1_writedata                (mm_interconnect_0_io_data_high_s1_writedata),               //                                   .writedata
		.io_data_high_s1_chipselect               (mm_interconnect_0_io_data_high_s1_chipselect),              //                                   .chipselect
		.io_data_low_s1_address                   (mm_interconnect_0_io_data_low_s1_address),                  //                     io_data_low_s1.address
		.io_data_low_s1_write                     (mm_interconnect_0_io_data_low_s1_write),                    //                                   .write
		.io_data_low_s1_readdata                  (mm_interconnect_0_io_data_low_s1_readdata),                 //                                   .readdata
		.io_data_low_s1_writedata                 (mm_interconnect_0_io_data_low_s1_writedata),                //                                   .writedata
		.io_data_low_s1_chipselect                (mm_interconnect_0_io_data_low_s1_chipselect),               //                                   .chipselect
		.io_riscv_flags_s1_address                (mm_interconnect_0_io_riscv_flags_s1_address),               //                  io_riscv_flags_s1.address
		.io_riscv_flags_s1_readdata               (mm_interconnect_0_io_riscv_flags_s1_readdata),              //                                   .readdata
		.jtag_uart_avalon_jtag_slave_address      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                   .write
		.jtag_uart_avalon_jtag_slave_read         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                   .read
		.jtag_uart_avalon_jtag_slave_readdata     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                   .chipselect
		.memory_s1_address                        (mm_interconnect_0_memory_s1_address),                       //                          memory_s1.address
		.memory_s1_write                          (mm_interconnect_0_memory_s1_write),                         //                                   .write
		.memory_s1_readdata                       (mm_interconnect_0_memory_s1_readdata),                      //                                   .readdata
		.memory_s1_writedata                      (mm_interconnect_0_memory_s1_writedata),                     //                                   .writedata
		.memory_s1_byteenable                     (mm_interconnect_0_memory_s1_byteenable),                    //                                   .byteenable
		.memory_s1_chipselect                     (mm_interconnect_0_memory_s1_chipselect),                    //                                   .chipselect
		.memory_s1_clken                          (mm_interconnect_0_memory_s1_clken),                         //                                   .clken
		.NiosII_debug_mem_slave_address           (mm_interconnect_0_niosii_debug_mem_slave_address),          //             NiosII_debug_mem_slave.address
		.NiosII_debug_mem_slave_write             (mm_interconnect_0_niosii_debug_mem_slave_write),            //                                   .write
		.NiosII_debug_mem_slave_read              (mm_interconnect_0_niosii_debug_mem_slave_read),             //                                   .read
		.NiosII_debug_mem_slave_readdata          (mm_interconnect_0_niosii_debug_mem_slave_readdata),         //                                   .readdata
		.NiosII_debug_mem_slave_writedata         (mm_interconnect_0_niosii_debug_mem_slave_writedata),        //                                   .writedata
		.NiosII_debug_mem_slave_byteenable        (mm_interconnect_0_niosii_debug_mem_slave_byteenable),       //                                   .byteenable
		.NiosII_debug_mem_slave_waitrequest       (mm_interconnect_0_niosii_debug_mem_slave_waitrequest),      //                                   .waitrequest
		.NiosII_debug_mem_slave_debugaccess       (mm_interconnect_0_niosii_debug_mem_slave_debugaccess)       //                                   .debugaccess
	);

	coprocessor_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (niosii_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (niosii_debug_reset_request_reset),   // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
